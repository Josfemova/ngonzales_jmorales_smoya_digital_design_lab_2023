module instr_rom
#(parameter WIDTH = 32, LENGTH = 1024)
(
	input clk, 
	input [(WIDTH-1):0] r_addr_a, r_addr_b,
	output logic [(WIDTH-1):0] rd_a, rd_b
);
	reg [(WIDTH-1):0] rom[(LENGTH-1):0];

	initial begin
		$readmemh("/home/josfemova/REPOSITORIOS/ngonzales_jmorales_smoya_digital_design_lab_2023/proyecto/rtl/memfile.dat",rom, 0, 22);
		//$readmemh("../code/build/program_le.txt", rom);
	end

	always @(posedge clk)
	begin
		rd_a <= rom[r_addr_a[WIDTH-1:2]];
		rd_b <= rom[r_addr_b[WIDTH-1:2]];
	end
endmodule
