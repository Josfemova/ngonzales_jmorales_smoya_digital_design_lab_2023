
module draw();

	
endmodule