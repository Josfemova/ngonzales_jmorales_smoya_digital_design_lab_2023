module laboratorio_3(
	input [3:0] A, B,	
	input [2:0] UC,
	output [3:0] Output,
	output [3:0] Flags	
);

endmodule