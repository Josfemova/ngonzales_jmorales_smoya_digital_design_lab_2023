package sprites;

parameter sprite_bg = 24'hf2e3c4;

const bit[23:0] color_bg = 24'hf2e3c4;
endpackage
